--
-- VHDL Architecture ece411.IR.untitled
--
-- Created:
--          by - page10.ews (linux6.ews.illinois.edu)
--          at - 20:25:51 01/21/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY IR IS
   PORT( 
      LoadIR       : IN     std_logic;
      MDRout       : IN     LC3b_word;
      SrcA         : OUT    LC3b_reg;
      SrcB         : OUT    LC3b_reg;
      imm5in       : OUT    LC3B_IMM5;
      offset9      : OUT    LC3b_offset9;
      opcode       : OUT    LC3b_opcode;
      clk          : IN     std_logic;
      imm5Flag     : OUT    std_logic;
      offset11Flag : OUT    std_logic;
      offset11     : OUT    LC3B_OFFSET11;
      IRDest       : OUT    LC3b_reg;
      index6       : OUT    LC3B_INDEX6;
      shiftType    : OUT    LC3B_SHFTOP;
      imm4in       : OUT    LC3B_SHIFTYPE;
      trapvect     : OUT    LC3B_TRAPVECT8
   );

-- Declarations

END IR ;

--
ARCHITECTURE UNTITLED OF IR IS
SIGNAL VAL_IR : LC3B_WORD;
BEGIN
	------------------------------
	VHDL_REG_IR : PROCESS (CLK, LOADIR, MDROUT)
	------------------------------
	BEGIN
		IF (CLK'EVENT AND (CLK = '1') AND (CLK'LAST_VALUE = '0')) THEN
			IF (LOADIR = '1') THEN
				VAL_IR <= MDROUT AFTER DELAY_REG;
			END IF;
		END IF;
	END PROCESS VHDL_REG_IR;
	OPCODE <= VAL_IR(15 DOWNTO 12);
	SRCA <= VAL_IR(8 DOWNTO 6);
	SRCB <= VAL_IR(2 DOWNTO 0);
	IRDest <= VAL_IR(11 DOWNTO 9);
	OFFSET9 <= VAL_IR(8 DOWNTO 0);
	imm5in <= VAL_IR(4 DOWNTO 0);
	INDEX6 <= VAL_IR(5 DOWNTO 0);
	imm5Flag<= VAL_IR(5);
	offset11Flag<=VAL_IR(11);
	offset11<=VAL_IR(10 DOWNTO 0);
	shiftType<=VAL_IR(5 downto 4);
	imm4in<=VAL_IR(3 downto 0);
	trapvect<=VAL_IR(7 downto 0);
END UNTITLED;

