--
-- VHDL Architecture ece411.ALU.untitled
--
-- Created:
--          by - page10.ews (linux6.ews.illinois.edu)
--          at - 20:22:46 01/21/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY ALU IS
   PORT( 
      ALUop     : IN     LC3b_aluop;
      RFAout    : IN     LC3b_word;
      ALUout    : OUT    LC3b_word;
      clk       : IN     std_logic;
      ALUMUXOUT : IN     LC3b_word
   );

-- Declarations

END ALU ;

--
ARCHITECTURE UNTITLED OF ALU IS
BEGIN
	----------------------------------------
	VHDL_ALU : PROCESS (RFAOUT, ALUMUXOUT, ALUOP)
	----------------------------------------
	VARIABLE TEMP_ALUOUT : LC3B_WORD;
	BEGIN
		-- CHECK FOR ALU OPERATION TYPE, AND EXECUTE
		CASE ALUOP IS
			WHEN ALU_ADD =>
				TEMP_ALUOUT := STD_LOGIC_VECTOR(SIGNED(RFAOUT) + SIGNED(ALUMUXOUT));
			WHEN ALU_AND =>
				TEMP_ALUOUT := (RFAOUT AND ALUMUXOUT);
			WHEN ALU_NOT =>
				TEMP_ALUOUT := (RFAOUT XOR "1111111111111111");
			WHEN ALU_PASS =>
				TEMP_ALUOUT := (RFAOUT);
			WHEN ALU_SLL=>
			  TEMP_ALUOUT := STD_LOGIC_VECTOR(SHIFT_LEFT(UNSIGNED(RFAOUT) , TO_INTEGER(UNSIGNED(ALUMUXOUT))));
			WHEN ALU_SRL=>
			  TEMP_ALUOUT := STD_LOGIC_VECTOR(SHIFT_RIGHT(UNSIGNED(RFAOUT) , TO_INTEGER(UNSIGNED(ALUMUXOUT))));
			WHEN ALU_SRA=>
			  TEMP_ALUOUT := STD_LOGIC_VECTOR(SHIFT_RIGHT(SIGNED(RFAOUT) , TO_INTEGER(UNSIGNED(ALUMUXOUT))));
			WHEN OTHERS =>
		END CASE;
	--SET OUTPUT VALUE ALUOUT TO BE THE TEMPORARY VALUE CALCULATED WITHIN THE PROCESS AFTER A DELAY
	ALUOUT <= TEMP_ALUOUT AFTER DELAY_ALU;
	END PROCESS VHDL_ALU;
END UNTITLED;
