--
-- VHDL Architecture ece411.Memory.untitled
--
-- Created:
--          by - page10.ews (linux6.ews.illinois.edu)
--          at - 21:30:53 01/21/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      Address   : IN     LC3b_word;
      DataOut   : IN     LC3B_WORD;
      MREAD_L   : IN     std_logic;
      MWRITEH_L : IN     std_logic;
      MWRITEL_L : IN     std_logic;
      RESET_L   : IN     std_logic;
      clk       : IN     std_logic;
      DataIn    : OUT    LC3B_WORD;
      MRESP_H   : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - page10.ews (gelib-057-02.ews.illinois.edu)
--          at - 14:57:33 03/01/13
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;


ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL ForceWrite   : std_logic;
   SIGNAL Miss         : std_logic;
   SIGNAL PMADDRESS    : LC3B_WORD;
   SIGNAL PMDATAIN     : LC3B_OWORD;
   SIGNAL PMDATAOUT    : LC3B_OWORD;
   SIGNAL PMREAD_L     : STD_LOGIC;
   SIGNAL PMRESP_H     : STD_LOGIC;
   SIGNAL PMWRITE_L    : STD_LOGIC;
   SIGNAL PickAddr     : STD_LOGIC;
   SIGNAL ReplaceCache : std_logic;
   SIGNAL WriteCache   : std_logic;
   SIGNAL dirtying     : std_logic;
   SIGNAL writeBack    : std_logic;


   -- Component Declarations
   COMPONENT Cache_Controller
   PORT (
      MREAD_L      : IN     std_logic ;
      Miss         : IN     std_logic ;
      PMRESP_H     : IN     STD_LOGIC ;
      RESET_L      : IN     std_logic ;
      ReplaceCache : IN     std_logic ;
      clk          : IN     std_logic ;
      dirtying     : IN     std_logic ;
      writeBack    : IN     std_logic ;
      ForceWrite   : OUT    std_logic ;
      PMREAD_L     : OUT    STD_LOGIC ;
      PMWRITE_L    : OUT    STD_LOGIC ;
      PickAddr     : OUT    STD_LOGIC ;
      WriteCache   : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Cache_Datapath
   PORT (
      Address      : IN     LC3b_word ;
      DataOut      : IN     LC3B_WORD ;
      ForceWrite   : IN     std_logic ;
      MREAD_L      : IN     std_logic ;
      MWRITEH_L    : IN     std_logic ;
      MWRITEL_L    : IN     std_logic ;
      PMDATAIN     : IN     LC3B_OWORD ;
      PickAddr     : IN     STD_LOGIC ;
      RESET_L      : IN     std_logic ;
      WriteCache   : IN     std_logic ;
      clk          : IN     std_logic ;
      DataIn       : OUT    LC3B_WORD ;
      Miss         : OUT    std_logic ;
      PMADDRESS    : OUT    LC3B_WORD ;
      PMDATAOUT    : OUT    LC3B_OWORD ;
      ReplaceCache : OUT    std_logic ;
      dirtying     : OUT    std_logic ;
      writeBack    : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Physical_Memory
   PORT (
      clk       : IN     std_logic ;
      PMADDRESS : IN     LC3B_WORD ;
      PMDATAOUT : IN     LC3B_OWORD ;
      PMREAD_L  : IN     STD_LOGIC ;
      RESET_L   : IN     std_logic ;
      PMDATAIN  : OUT    LC3B_OWORD ;
      PMRESP_H  : OUT    STD_LOGIC ;
      PMWRITE_L : IN     STD_LOGIC 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Controller USE ENTITY ece411.Cache_Controller;
   FOR ALL : Cache_Datapath USE ENTITY ece411.Cache_Datapath;
   FOR ALL : Physical_Memory USE ENTITY ece411.Physical_Memory;
   -- pragma synthesis_on


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 eb1
   -- eb1 1 
   MRESP_H<=not(miss);                                       


   -- Instance port mappings.
   Cache_Cont : Cache_Controller
      PORT MAP (
         MREAD_L      => MREAD_L,
         Miss         => Miss,
         PMRESP_H     => PMRESP_H,
         RESET_L      => RESET_L,
         ReplaceCache => ReplaceCache,
         clk          => clk,
         dirtying     => dirtying,
         writeBack    => writeBack,
         ForceWrite   => ForceWrite,
         PMREAD_L     => PMREAD_L,
         PMWRITE_L    => PMWRITE_L,
         PickAddr     => PickAddr,
         WriteCache   => WriteCache
      );
   Cache_DP : Cache_Datapath
      PORT MAP (
         Address      => Address,
         DataOut      => DataOut,
         ForceWrite   => ForceWrite,
         MREAD_L      => MREAD_L,
         MWRITEH_L    => MWRITEH_L,
         MWRITEL_L    => MWRITEL_L,
         PMDATAIN     => PMDATAIN,
         PickAddr     => PickAddr,
         RESET_L      => RESET_L,
         WriteCache   => WriteCache,
         clk          => clk,
         DataIn       => DataIn,
         Miss         => Miss,
         PMADDRESS    => PMADDRESS,
         PMDATAOUT    => PMDATAOUT,
         ReplaceCache => ReplaceCache,
         dirtying     => dirtying,
         writeBack    => writeBack
      );
   PDRAM : Physical_Memory
      PORT MAP (
         clk       => clk,
         PMADDRESS => PMADDRESS,
         PMDATAOUT => PMDATAOUT,
         PMREAD_L  => PMREAD_L,
         RESET_L   => RESET_L,
         PMDATAIN  => PMDATAIN,
         PMRESP_H  => PMRESP_H,
         PMWRITE_L => PMWRITE_L
      );

END struct;
